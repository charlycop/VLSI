* polarisation d'un transistor NMOS


* La commande .INCLUDE permet d'inserer le contenu d'un fichier
.include ../mosn_mosp.wc

* instanciation du transistor NMOS
MN dd grille 0 0 TN L=0.35e-06 W=1.4e-06

* declaration des source de tensions
Vd dd 0 dc 3.3
Vg grille 0 dc 3.3

* Analyse statique
.DC Vg 0.0 3.3 {3.3/63}
*.DC Vd 0.0 3.3 {3.3/63} vg 0 3.3 0.5

* affichage des resultats
.PLOT ID(MN)

* fin de la description du circuit 
.END

* Spice description of buf_x8
* Spice driver version 1169777
* Date ( dd/mm/yyyy hh:mm:ss ):  5/10/2006 at 14:32:30

* INTERF i q vdd vss 

.lib typical
.include ../mosn_mosp.wc
.lib "buf_x8.spi" circuit
.endl  typical

.lib circuit

.subckt buf_x8 2 52 16 41 
* NET 2 = i
* NET 16 = vdd
* NET 41 = vss
* NET 52 = q
Mtr_00010 56 33 6 16 tp L=0.35U W=5.9U AS=4.425P AD=4.425P PS=13.3U PD=13.3U 
Mtr_00009 7 34 56 16 tp L=0.35U W=5.9U AS=4.425P AD=4.425P PS=13.3U PD=13.3U 
Mtr_00008 57 35 7 16 tp L=0.35U W=5.9U AS=4.425P AD=4.425P PS=13.3U PD=13.3U 
Mtr_00007 9 36 57 16 tp L=0.35U W=5.9U AS=4.425P AD=4.425P PS=13.3U PD=13.3U 
Mtr_00006 6 3 31 16 tp L=0.35U W=5.9U AS=4.425P AD=4.425P PS=13.3U PD=13.3U 
Mtr_00005 51 22 43 41 tn L=0.35U W=2.9U AS=2.175P AD=2.175P PS=7.3U PD=7.3U 
Mtr_00004 42 21 51 41 tn L=0.35U W=2.9U AS=2.175P AD=2.175P PS=7.3U PD=7.3U 
Mtr_00003 43 23 53 41 tn L=0.35U W=2.9U AS=2.175P AD=2.175P PS=7.3U PD=7.3U 
Mtr_00002 53 24 44 41 tn L=0.35U W=2.9U AS=2.175P AD=2.175P PS=7.3U PD=7.3U 
Mtr_00001 19 1 42 41 tn L=0.35U W=2.9U AS=2.175P AD=2.175P PS=7.3U PD=7.3U 
R5_1 1 2 12
R5_2 3 2 12
R4_1 6 16 12
R4_2 9 16 12
R4_3 7 16 12
R4_4 9 15 12
R4_5 7 8 12
R4_6 7 11 12
R4_7 7 14 12
R4_8 10 13 0.087
C4_81 10 41 1.46887e-16
C4_82 13 41 1.46887e-16
R4_9 12 13 0.087
C4_91 12 41 1.1751e-16
C4_92 13 41 1.1751e-16
R4_10 14 16 0.174
C4_101 14 41 2.05643e-16
C4_102 16 41 2.05643e-16
R4_11 11 14 0.087
C4_111 11 41 1.46887e-16
C4_112 14 41 1.46887e-16
R4_12 8 11 0.087
C4_121 8 41 1.46887e-16
C4_122 11 41 1.46887e-16
R4_13 15 16 0.174
C4_131 15 41 2.05643e-16
C4_132 16 41 2.05643e-16
R4_14 12 15 0.174
C4_141 12 41 1.76265e-16
C4_142 15 41 1.76265e-16
R3_1 19 20 12
R3_2 31 32 12
R3_3 31 37 12
R3_4 31 38 12
R3_5 26 25 12
R3_6 27 33 90
C3_61 27 41 6.07294e-16
C3_62 33 41 6.07294e-16
R3_7 21 27 60
C3_71 21 41 4.33781e-16
C3_72 27 41 4.33781e-16
R3_8 29 35 90
C3_81 29 41 6.07294e-16
C3_82 35 41 6.07294e-16
R3_9 23 29 60
C3_91 23 41 4.33781e-16
C3_92 29 41 4.33781e-16
R3_10 28 34 90
C3_101 28 41 6.07294e-16
C3_102 34 41 6.07294e-16
R3_11 22 28 60
C3_111 22 41 4.33781e-16
C3_112 28 41 4.33781e-16
R3_12 30 36 90
C3_121 30 41 6.07294e-16
C3_122 36 41 6.07294e-16
R3_13 24 30 60
C3_131 24 41 4.33781e-16
C3_132 30 41 4.33781e-16
R3_14 29 30 6
C3_141 29 41 2.62755e-16
C3_142 30 41 2.62755e-16
R3_15 28 29 6
C3_151 28 41 2.62755e-16
C3_152 29 41 2.62755e-16
R3_16 27 28 6
C3_161 27 41 2.62755e-16
C3_162 28 41 2.62755e-16
R3_17 26 27 12
C3_171 26 41 3.94133e-16
C3_172 27 41 3.94133e-16
R3_18 38 37 0.174
C3_181 38 41 1.40925e-16
C3_182 37 41 1.40925e-16
R3_19 32 38 0.174
C3_191 32 41 1.40925e-16
C3_192 38 41 1.40925e-16
R3_20 25 32 0.435
C3_201 25 41 2.8185e-16
C3_202 32 41 2.8185e-16
R3_21 20 25 0.435
C3_211 20 41 2.8185e-16
C3_212 25 41 2.8185e-16
R2_1 43 41 12
R2_2 43 45 12
R2_3 44 41 12
R2_4 42 41 12
R2_5 44 46 12
R2_6 47 48 0.087
C2_61 47 41 1.1751e-16
C2_62 48 41 1.1751e-16
R2_7 46 47 0.174
C2_71 46 41 2.05643e-16
C2_72 47 41 2.05643e-16
R2_8 41 46 0.174
C2_81 41 41 2.05643e-16
C2_82 46 41 2.05643e-16
R2_9 41 45 0.174
C2_91 41 41 2.05643e-16
C2_92 45 41 2.05643e-16
R1_1 51 52 12
R1_2 56 52 4
R1_3 59 57 12
R1_4 60 57 12
R1_5 58 57 12
R1_6 54 53 12
R1_7 59 60 0.087
C1_71 59 41 1.46887e-16
C1_72 60 41 1.46887e-16
R1_8 58 59 0.087
C1_81 58 41 1.46887e-16
C1_82 59 41 1.46887e-16
R1_9 55 58 0.261
C1_91 55 41 2.93775e-16
C1_92 58 41 2.93775e-16
R1_10 54 55 0.261
C1_101 54 41 2.93775e-16
C1_102 55 41 2.93775e-16
R1_11 52 55 0.348
C1_111 52 41 3.5253e-16
C1_112 55 41 3.5253e-16
.ends buf_x8
.endl circuit
